magic
tech sky130A
magscale 1 2
timestamp 1597433933
<< error_p >>
rect -109 6 109 42
rect -109 -78 -73 6
rect 73 -78 109 6
rect -109 -114 109 -78
<< pmos >>
rect -15 -78 15 6
<< pdiff >>
rect -73 -6 -15 6
rect -73 -66 -61 -6
rect -27 -66 -15 -6
rect -73 -78 -15 -66
rect 15 -6 73 6
rect 15 -66 27 -6
rect 61 -66 73 -6
rect 15 -78 73 -66
<< pdiffc >>
rect -61 -66 -27 -6
rect 27 -66 61 -6
<< poly >>
rect -33 87 33 103
rect -33 53 -17 87
rect 17 53 33 87
rect -33 37 33 53
rect -15 6 15 37
rect -15 -104 15 -78
<< polycont >>
rect -17 53 17 87
<< locali >>
rect -33 53 -17 87
rect 17 53 33 87
rect -61 -6 -27 10
rect -61 -82 -27 -66
rect 27 -6 61 10
rect 27 -82 61 -66
<< properties >>
string gencell pshort
string parameters w 0.42 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {pshort plowvt phighvt phv} full_metal 1
string library sky130
<< end >>
