magic
tech sky130A
magscale 1 2
timestamp 1597433202
<< nwell >>
rect -163 -80 164 89
<< pmos >>
rect -63 -42 -33 42
rect 33 -42 63 42
<< pdiff >>
rect -125 30 -63 42
rect -125 -30 -113 30
rect -79 -30 -63 30
rect -125 -42 -63 -30
rect -33 30 33 42
rect -33 -30 -17 30
rect 17 -30 33 30
rect -33 -42 33 -30
rect 63 30 125 42
rect 63 -30 79 30
rect 113 -30 125 30
rect 63 -42 125 -30
<< pdiffc >>
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
<< poly >>
rect -63 42 -33 68
rect 33 42 63 68
rect -63 -73 -33 -42
rect 33 -73 63 -42
rect -81 -139 81 -73
<< locali >>
rect -113 30 -79 46
rect -113 -46 -79 -30
rect -17 30 17 46
rect -17 -46 17 -30
rect 79 30 113 46
rect 79 -46 113 -30
<< labels >>
rlabel pdiffc -17 -30 17 30 1 Vdd!
rlabel pdiffc -113 -30 -79 30 1 Vout_pos
rlabel pdiffc 79 -30 113 30 1 Vout_neg
rlabel poly -81 -139 81 -73 1 Vbias2
<< properties >>
string gencell pshort
string parameters w 0.42 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {pshort plowvt phighvt phv} full_metal 1
string library sky130
<< end >>
